//===========================================================================
// Module name: key_test.v
// Описание: Обнаружьте 2 кнопки KEY1 ~ KEY2 на плате разработки, когда кнопка обнаружена, светодиодный индикатор перевернется
//===========================================================================
`timescale 1ns / 1ps
module key_test  (
							clk,              // Входные часы на плате разработки: 50Mhz
							rst_n,            // вводим кнопку сброса на отладочной плате
							key_in,           // Ввод сигнала ключа (KEY1 ~ KEY2)
							led_out           // Выход, используемый для управления светодиодом на плате разработки
						);

//===========================================================================
// PORT declarations
//===========================================================================						
input        clk; 
input        rst_n;
input  [1:0] key_in;
output 		 led_out;

//Определение регистра
reg [19:0] count;
reg [1:0] key_scan; //Значение сканирования ключа KEY

//===========================================================================
// Выборка значения кнопки, сканирование один раз в 20 мс, частота выборки меньше, чем частота сбоев кнопки, что эквивалентно фильтрации высокочастотного сигнала сбоя.
//===========================================================================
always @(posedge clk or negedge rst_n)     //Обнаружение нарастающего фронта часов и спадающего фронта сброса
begin
   if(!rst_n)                //Активный сигнал сброса низкий
      count <= 20'd0;        //Счетчик очищен
   else
      begin
         if(count ==20'd999_999)   //Сканируйте кнопку за 20 мс, считайте за 20 мс (50M / 50-1 = 999_999)
            begin
               count <= 20'b0;     //Счетчик считает до 20 мс, и счетчик очищается.
               key_scan <= key_in; //Уровень входного сигнала сэмплирования
            end
         else
            count <= count + 20'b1; //Счетчик плюс 1
     end
end
//===========================================================================
// Сигнал ключа фиксирует такт часов
//===========================================================================
reg [1:0] key_scan_r;
always @(posedge clk)
    key_scan_r <= key_scan;       
    
wire [1:0] flag_key = key_scan_r[1:0] & (~key_scan[1:0]);  //Когда обнаруживается изменение спадающего фронта кнопки, это означает, что кнопка нажата и кнопка действительна.

//===========================================================================
// Управление светодиодной подсветкой, когда кнопка нажата, соответствующий светодиодный выход меняется на противоположный
//===========================================================================
reg temp_led;
always @ (posedge clk or negedge rst_n)      //Обнаружение нарастающего фронта часов и спадающего фронта сброса
begin
    if (!rst_n)                 					//Активный сигнал сброса низкий
         temp_led <= 1'b1;   						//Выходной сигнал управления светодиодной подсветкой низкий, светодиодная подсветка не горит
    else
         begin            
             if ( flag_key[0] ) temp_led <= ~temp_led;   //При изменении значения KEY1 светодиод будет включаться и выключаться.
             if ( flag_key[1] ) temp_led <= ~temp_led;   //При изменении значения KEY2 светодиод будет включаться и выключаться.
         end
end
 
 assign led_out = temp_led;

endmodule

