/***************************************/
// Модуль кодирования: десятичное число -> 7-сегментная цифровая трубка       //
/***************************************/
module smg_encode_module
(
	 input CLK,
	 input RSTn,
	 input [3:0]Number_Data,
	 output [6:0]SMG_Data
);

	 /***************************************/
	 
	 parameter _0 = 7'b100_0000, _1 = 7'b111_1001, _2 = 7'b010_0100, 
	           _3 = 7'b011_0000, _4 = 7'b001_1001, _5 = 7'b001_0010, 
				  _6 = 7'b000_0010, _7 = 7'b111_1000, _8 = 7'b000_0000,
				  _9 = 7'b001_0000;
	 
	 /***************************************/
	 
	 reg [6:0]rSMG;

	 always @ ( posedge CLK or negedge RSTn )
	     if( !RSTn )
		      begin
				    rSMG <= 7'b111_1111;
				end
        else 
		       case( Number_Data )
		           
					  4'd0 : rSMG <= _0;
					  4'd1 : rSMG <= _1;
					  4'd2 : rSMG <= _2;
					  4'd3 : rSMG <= _3;
					  4'd4 : rSMG <= _4;
					  4'd5 : rSMG <= _5;
					  4'd6 : rSMG <= _6;
					  4'd7 : rSMG <= _7;
					  4'd8 : rSMG <= _8;
					  4'd9 : rSMG <= _9;
					  
				 endcase
		      
	 /***************************************/
	 
	 assign SMG_Data = rSMG;
	 
	 /***************************************/
			  
endmodule
