`timescale 1ns / 1ps

module led_test (
                  clk,           // Входные часы на плате разработки: 50Mhz
                  rst_n,         // вводим кнопку сброса на отладочной плате
                  led            // выходной светодиодный индикатор
             );
             
//===========================================================================
// PORT declarations
//===========================================================================
input clk;
input rst_n;
output led;

//Определение регистра
reg [31:0] timer;                  
reg led;


//===========================================================================
// Счетчик счетчика: счетчик циклов 0 ~ 2 секунды
//===========================================================================
  always @(posedge clk or negedge rst_n)    //Обнаружение нарастающего фронта часов и спадающего фронта сброса
    begin
      if (~rst_n)                           //Активный сигнал сброса низкий
          timer <= 0;                       //Сброс счетчика
      else if (timer == 32'd99_999_999)     //Кварцевый генератор, используемый платой разработки, составляет 50 МГц, счетчик 2 секунды (50M*2-1=99_999_999)
          timer <= 0;                       //Счетчик считает до 2 секунд, счетчик обнуляется.
      else
		    timer <= timer + 1'b1;            //Счетчик плюс 1
    end

//===========================================================================
// LED Контроль света
//===========================================================================
  always @(posedge clk or negedge rst_n)   //Обнаружение нарастающего фронта часов и спадающего фронта сброса
    begin
      if (~rst_n)                          //Активный сигнал сброса низкий
          led <= 1'b1;                  	 //LED 
      else if (timer == 32'd49_999_999)    //Счетчик считает до 1 секунды,
          led <= 1'b0;                     //LED Загораться
      else if (timer == 32'd99_999_999)    //Счетчик считает до 2 секунд,
          led <= 1'b1;                     //LED Гаснет
    end
endmodule

