library verilog;
use verilog.vl_types.all;
entity pll_test_tb is
end pll_test_tb;
