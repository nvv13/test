module test1_bl



endmodule

